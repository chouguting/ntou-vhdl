library verilog;
use verilog.vl_types.all;
entity generic_multiplier_8bit_vlg_vec_tst is
end generic_multiplier_8bit_vlg_vec_tst;
