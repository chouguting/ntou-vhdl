library verilog;
use verilog.vl_types.all;
entity counter_20_to_A0_vlg_vec_tst is
end counter_20_to_A0_vlg_vec_tst;
