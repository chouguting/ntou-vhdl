library verilog;
use verilog.vl_types.all;
entity generic_shift_register_8bit_ex_vlg_vec_tst is
end generic_shift_register_8bit_ex_vlg_vec_tst;
