library verilog;
use verilog.vl_types.all;
entity bcd_counter_100_to_499_vlg_vec_tst is
end bcd_counter_100_to_499_vlg_vec_tst;
