library verilog;
use verilog.vl_types.all;
entity clk_with_number_vlg_vec_tst is
end clk_with_number_vlg_vec_tst;
