library verilog;
use verilog.vl_types.all;
entity BCD_cascading_counter_12bit_vlg_vec_tst is
end BCD_cascading_counter_12bit_vlg_vec_tst;
