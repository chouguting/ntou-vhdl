library verilog;
use verilog.vl_types.all;
entity div_20 is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        P               : out    vl_logic
    );
end div_20;
