library verilog;
use verilog.vl_types.all;
entity adder_subtractor_arithmetic_vlg_vec_tst is
end adder_subtractor_arithmetic_vlg_vec_tst;
