library verilog;
use verilog.vl_types.all;
entity clk_count_0000_to_9999_vlg_vec_tst is
end clk_count_0000_to_9999_vlg_vec_tst;
