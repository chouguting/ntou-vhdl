library verilog;
use verilog.vl_types.all;
entity mux8_1_vlg_check_tst is
    port(
        D_out           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux8_1_vlg_check_tst;
