library verilog;
use verilog.vl_types.all;
entity adder_14bits_vlg_vec_tst is
end adder_14bits_vlg_vec_tst;
