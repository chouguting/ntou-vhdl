library verilog;
use verilog.vl_types.all;
entity step_wave_vlg_vec_tst is
end step_wave_vlg_vec_tst;
