library verilog;
use verilog.vl_types.all;
entity adder_1bit_vlg_vec_tst is
end adder_1bit_vlg_vec_tst;
