library verilog;
use verilog.vl_types.all;
entity breathing_light_5sec_vlg_vec_tst is
end breathing_light_5sec_vlg_vec_tst;
