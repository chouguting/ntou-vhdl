library verilog;
use verilog.vl_types.all;
entity generate_demux_1to8_vlg_vec_tst is
end generate_demux_1to8_vlg_vec_tst;
