library verilog;
use verilog.vl_types.all;
entity fast_multiplier_8bit_vlg_vec_tst is
end fast_multiplier_8bit_vlg_vec_tst;
