library verilog;
use verilog.vl_types.all;
entity div_20_vlg_check_tst is
    port(
        P               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end div_20_vlg_check_tst;
