library verilog;
use verilog.vl_types.all;
entity mux8_1_vlg_vec_tst is
end mux8_1_vlg_vec_tst;
