library verilog;
use verilog.vl_types.all;
entity generic_adder_8bit_vlg_vec_tst is
end generic_adder_8bit_vlg_vec_tst;
